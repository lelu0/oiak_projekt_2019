//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "pic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w6;    //: /sn:0 {0}(157,415)(139,415){1}
//: {2}(135,415)(111,415)(111,396)(98,396){3}
//: {4}(137,417)(137,487)(206,487){5}
reg w4;    //: /sn:0 {0}(607,279)(663,279)(663,238)(677,238){1}
reg [7:0] w0;    //: /sn:0 {0}(#:108,264)(108,274)(239,274)(239,284){1}
//: {2}(241,286)(247,286){3}
//: {4}(237,286)(#:230,286){5}
reg w3;    //: /sn:0 {0}(606,194)(662,194)(662,233)(677,233){1}
reg [7:0] w1;    //: /sn:0 {0}(#:105,357)(105,367)(243,367)(243,320){1}
//: {2}(245,318)(247,318){3}
//: {4}(241,318)(#:230,318){5}
reg w8;    //: /sn:0 {0}(157,420)(119,420)(119,446)(113,446){1}
//: {2}(109,446)(98,446){3}
//: {4}(111,448)(111,492)(206,492){5}
reg w10;    //: /sn:0 {0}(100,494)(124,494)(124,446)(192,446)(192,441){1}
//: {2}(194,439)(201,439)(201,456)(207,456){3}
//: {4}(192,437)(192,423)(214,423){5}
reg w5;    //: /sn:0 {0}(261,278)(261,253)(285,253){1}
wire [7:0] w7;    //: /sn:0 {0}(#:276,302)(283,302){1}
//: {2}(287,302)(293,302){3}
//: {4}(285,300)(#:285,290)(399,290)(399,268){5}
wire w14;    //: /sn:0 {0}(277,401)(277,421)(235,421){1}
wire w16;    //: /sn:0 {0}(228,459)(250,459)(250,470)(265,470){1}
wire w19;    //: /sn:0 {0}(227,490)(250,490)(250,475)(265,475){1}
wire w15;    //: /sn:0 {0}(320,454)(320,473)(286,473){1}
wire w2;    //: /sn:0 {0}(698,236)(757,236)(757,214){1}
wire w13;    //: /sn:0 {0}(214,418)(201,418)(201,418)(186,418){1}
//: {2}(184,416)(184,461)(207,461){3}
//: {4}(182,418)(178,418){5}
wire w9;    //: /sn:0 {0}(261,326)(261,341){1}
//: enddecls

  //: joint g8 (w1) @(243, 318) /w:[ 2 -1 4 1 ]
  //: DIP g4 (w0) @(108,254) /sn:0 /w:[ 0 ] /st:3 /dn:1
  //: SWITCH g3 (w4) @(590,279) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g13 (w8) @(81,446) /sn:0 /w:[ 3 ] /st:1 /dn:1
  //: SWITCH g2 (w3) @(589,194) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g1 (w2) @(757,207) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g11 (w5) @(303,253) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  _GGXOR2 #(8) g16 (.I0(w13), .I1(w10), .Z(w14));   //: @(225,421) /sn:0 /w:[ 0 5 1 ]
  //: joint g10 (w7) @(285, 302) /w:[ 2 4 1 -1 ]
  //: joint g19 (w10) @(192, 439) /w:[ 2 4 -1 1 ]
  _GGADD8 #(68, 70, 62, 64) g6 (.A(w1), .B(w0), .S(w7), .CI(w5), .CO(w9));   //: @(263,302) /sn:0 /R:1 /w:[ 3 3 0 0 0 ]
  //: LED g9 (w7) @(399,261) /sn:0 /w:[ 5 ] /type:1
  //: joint g7 (w0) @(239, 286) /w:[ 2 1 4 -1 ]
  _GGXOR2 #(8) g15 (.I0(w6), .I1(w8), .Z(w13));   //: @(168,418) /sn:0 /w:[ 0 0 5 ]
  //: joint g20 (w13) @(184, 418) /w:[ 1 2 4 -1 ]
  _GGAND2 #(6) g17 (.I0(w10), .I1(w13), .Z(w16));   //: @(218,459) /sn:0 /w:[ 3 3 0 ]
  //: LED g25 (w15) @(320,447) /sn:0 /w:[ 0 ] /type:0
  //: DIP g5 (w1) @(105,347) /sn:0 /w:[ 0 ] /st:3 /dn:1
  //: SWITCH g14 (w10) @(83,494) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g21 (w8) @(111, 446) /w:[ 1 -1 2 4 ]
  //: LED g24 (w14) @(277,394) /sn:0 /w:[ 0 ] /type:0
  _GGOR2 #(6) g23 (.I0(w16), .I1(w19), .Z(w15));   //: @(276,473) /sn:0 /w:[ 1 1 1 ]
  _GGAND2 #(6) g0 (.I0(w3), .I1(w4), .Z(w2));   //: @(688,236) /sn:0 /w:[ 1 1 0 ]
  //: joint g22 (w6) @(137, 415) /w:[ 1 -1 2 4 ]
  //: SWITCH g12 (w6) @(81,396) /sn:0 /w:[ 3 ] /st:0 /dn:1
  _GGAND2 #(6) g18 (.I0(w6), .I1(w8), .Z(w19));   //: @(217,490) /sn:0 /w:[ 5 5 0 ]

endmodule
//: /netlistEnd

