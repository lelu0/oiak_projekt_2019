//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w4;    //: /sn:0 {0}(607,279)(663,279)(663,238)(677,238){1}
reg [7:0] w0;    //: /sn:0 {0}(#:78,197)(78,207)(209,207)(209,217){1}
//: {2}(211,219)(217,219){3}
//: {4}(207,219)(#:200,219){5}
reg w3;    //: /sn:0 {0}(606,194)(662,194)(662,233)(677,233){1}
reg [7:0] w1;    //: /sn:0 {0}(#:75,290)(75,300)(213,300)(213,253){1}
//: {2}(215,251)(217,251){3}
//: {4}(211,251)(#:200,251){5}
reg w5;    //: /sn:0 {0}(231,211)(231,136)(254,136){1}
wire [7:0] w7;    //: /sn:0 {0}(#:246,235)(253,235){1}
//: {2}(257,235)(263,235){3}
//: {4}(255,233)(#:255,223)(369,223)(369,201){5}
wire w2;    //: /sn:0 {0}(698,236)(757,236)(757,214){1}
wire w9;    //: /sn:0 {0}(231,259)(231,274){1}
//: enddecls

  //: joint g8 (w1) @(213, 251) /w:[ 2 -1 4 1 ]
  //: DIP g4 (w0) @(78,187) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g3 (w4) @(590,279) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: SWITCH g2 (w3) @(589,194) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g1 (w2) @(757,207) /sn:0 /w:[ 1 ] /type:0
  //: SWITCH g11 (w5) @(272,136) /sn:0 /R:2 /w:[ 1 ] /st:0 /dn:1
  //: joint g10 (w7) @(255, 235) /w:[ 2 4 1 -1 ]
  _GGADD8 #(68, 70, 62, 64) g6 (.A(w1), .B(w0), .S(w7), .CI(w5), .CO(w9));   //: @(233,235) /sn:0 /R:1 /w:[ 3 3 0 0 0 ]
  //: LED g9 (w7) @(369,194) /sn:0 /w:[ 5 ] /type:1
  //: joint g7 (w0) @(209, 219) /w:[ 2 1 4 -1 ]
  //: DIP g5 (w1) @(75,280) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGAND2 #(6) g0 (.I0(w3), .I1(w4), .Z(w2));   //: @(688,236) /sn:0 /w:[ 1 1 0 ]

endmodule
//: /netlistEnd

