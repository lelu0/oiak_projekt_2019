//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "pic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg w1;    //: /sn:0 {0}(229,160)(235,160)(235,120){1}
supply1 w8;    //: /sn:0 {0}(389,160)(479,160)(479,133){1}
supply0 w11;    //: /sn:0 {0}(507,182)(399,182)(399,170)(389,170){1}
supply1 w5;    //: /sn:0 {0}(54,109)(54,151)(66,151)(66,160){1}
reg [7:0] w9;    //: /sn:0 {0}(#:276,299)(276,284){1}
wire w6;    //: /sn:0 {0}(285,203)(305,203)(305,194){1}
//: {2}(305,190)(305,165)(313,165){3}
//: {4}(303,192)(288,192)(288,182)(229,182)(229,246)(71,246)(71,236){5}
wire [11:0] w7;    //: /sn:0 {0}(#:357,83)(357,93)(350,93){1}
//: {2}(349,93)(#:252,93){3}
wire w14;    //: /sn:0 {0}(198,311)(183,311){1}
wire [9:0] w4;    //: /sn:0 {0}(#:81,198)(125,198){1}
//: {2}(#:129,198)(143,198)(143,297){3}
//: {4}(127,196)(127,131){5}
//: {6}(129,129)(139,129)(139,95)(#:217,95){7}
//: {8}(127,127)(127,121){9}
wire w15;    //: /sn:0 {0}(135,311)(120,311){1}
wire [9:0] w0;    //: /sn:0 {0}(#:159,326)(159,397)(106,397){1}
//: {2}(#:102,397)(75,397)(75,320){3}
//: {4}(104,399)(104,431)(#:18,431)(18,198)(60,198){5}
wire [5:0] w3;    //: /sn:0 {0}(#:350,97)(350,155){1}
wire [5:0] w2;    //: /sn:0 {0}(#:350,176)(350,191){1}
wire [9:0] w12;    //: /sn:0 {0}(#:275,285)(175,285)(175,297){1}
wire w10;    //: /sn:0 {0}(71,48)(98,48)(98,138)(76,138)(76,160){1}
//: enddecls

  //: VDD g4 (w8) @(490,133) /sn:0 /w:[ 1 ]
  _GGREG10 #(10, 10, 20) g8 (.Q(w4), .D(w0), .EN(w10), .CLR(w5), .CK(w6));   //: @(71,198) /sn:0 /R:1 /w:[ 0 5 1 1 5 ]
  _GGREG6 #(10, 10, 20) g3 (.Q(w2), .D(w3), .EN(w11), .CLR(w8), .CK(w6));   //: @(350,165) /sn:0 /w:[ 0 1 1 0 3 ]
  _GGCLOCK_P3000_0_50 g13 (.Z(w10));   //: @(58,48) /sn:0 /w:[ 0 ] /omega:3000 /phi:0 /duty:50
  //: SWITCH g2 (w1) @(212,160) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g1 (w4) @(127, 198) /w:[ 2 4 1 -1 ]
  //: joint g11 (w6) @(305, 192) /w:[ -1 2 4 1 ]
  //: comment g16 @(355,139) /sn:0
  //: /line:"Instruction register"
  //: /line:""
  //: /end
  //: joint g10 (w4) @(127, 129) /w:[ 6 8 -1 5 ]
  //: LED g19 (w0) @(75,313) /sn:0 /w:[ 3 ] /type:1
  _GGCLOCK_P100_0_50 g6 (.Z(w6));   //: @(272,203) /sn:0 /w:[ 0 ] /omega:100 /phi:0 /duty:50
  assign w3 = w7[5:0]; //: TAP g7 @(350,91) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: LED g9 (w7) @(357,76) /sn:0 /w:[ 0 ] /type:1
  //: joint g20 (w0) @(104, 397) /w:[ 1 -1 2 4 ]
  //: comment g15 @(192,52) /sn:0
  //: /line:"Program memory"
  //: /end
  _GGADD10 #(84, 86, 78, 80) g17 (.A(w4), .B(w12), .S(w0), .CI(w14), .CO(w15));   //: @(159,313) /sn:0 /w:[ 3 1 0 1 0 ]
  //: comment g14 @(85,206) /sn:0
  //: /line:"Program counter"
  //: /line:""
  //: /end
  //: GROUND g5 (w11) @(513,182) /sn:0 /R:1 /w:[ 0 ]
  _GGROM10x12 #(10, 30) g0 (.A(w4), .D(w7), .OE(w1));   //: @(235,94) /sn:0 /w:[ 7 3 1 ] /mem:"/home/lelu0/oiakp/program.mem"
  //: VDD g12 (w5) @(65,109) /sn:0 /w:[ 0 ]
  //: DIP g18 (w9) @(276,310) /sn:0 /R:2 /w:[ 0 ] /st:1 /dn:1

endmodule
//: /netlistEnd

//: /netlistBegin ROM
module ROM();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
reg [7:0] w1;    //: /sn:0 {0}(#:92,155)(92,159){1}
//: {2}(94,161)(#:104,161)(104,250)(169,250){3}
//: {4}(92,163)(92,172){5}
reg w2;    //: /sn:0 {0}(121,324)(175,324)(175,282)(185,282){1}
//: {2}(187,280)(187,275){3}
//: {4}(187,284)(187,292){5}
wire [7:0] w0;    //: /sn:0 {0}(#:204,248)(267,248)(267,166)(277,166){1}
//: {2}(279,164)(279,158){3}
//: {4}(279,168)(#:279,175){5}
//: enddecls

  //: joint g4 (w0) @(279, 166) /w:[ -1 2 1 4 ]
  //: joint g3 (w1) @(92, 161) /w:[ 2 1 -1 4 ]
  _GGROM8x8 #(10, 30) g2 (.A(w1), .D(w0), .OE(w2));   //: @(187,249) /sn:0 /w:[ 3 0 3 ]
  //: DIP g1 (w1) @(92,145) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g6 (w2) @(187, 282) /w:[ -1 2 1 4 ]
  //: SWITCH g5 (w2) @(104,324) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g0 (w0) @(279,151) /sn:0 /w:[ 3 ] /type:1

endmodule
//: /netlistEnd

