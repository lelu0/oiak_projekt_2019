//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "pic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
supply0 w16;    //: /sn:0 {0}(206,330)(206,311)(183,311){1}
supply1 w15;    //: /sn:0 {0}(734,224)(734,253)(715,253)(715,238){1}
reg w0;    //: /sn:0 {0}(46,48)(96,48){1}
//: {2}(100,48)(130,48)(130,22){3}
//: {4}(98,50)(98,142)(75,142)(75,160){5}
reg w1;    //: /sn:0 {0}(229,160)(235,160)(235,120){1}
supply1 w8;    //: /sn:0 {0}(389,160)(445,160)(445,157){1}
//: {2}(447,155)(477,155)(477,47)(544,47)(544,57){3}
//: {4}(445,153)(445,135){5}
supply0 w18;    //: /sn:0 {0}(689,302)(689,315){1}
//: {2}(691,317)(705,317)(705,238){3}
//: {4}(689,319)(689,510)(674,510){5}
supply0 w11;    //: /sn:0 {0}(439,91)(422,91){1}
//: {2}(418,91)(402,91)(402,168){3}
//: {4}(404,170)(420,170)(420,439)(465,439)(465,429){5}
//: {6}(400,170)(389,170){7}
//: {8}(420,93)(420,121)(535,121){9}
//: {10}(539,121)(551,121)(551,107){11}
//: {12}(537,119)(537,107){13}
reg [7:0] w10;    //: /sn:0 {0}(#:882,627)(882,637)(758,637)(758,343){1}
reg w13;    //: /sn:0 {0}(47,94)(65,94)(65,160){1}
reg [8:0] w9;    //: /sn:0 {0}(#:317,361)(317,290)(177,290){1}
//: {2}(175,288)(#:175,283){3}
//: {4}(175,292)(175,297){5}
wire w6;    //: /sn:0 {0}(379,469)(372,469)(372,471)(347,471){1}
wire [7:0] acc_in;    //: /sn:0 {0}(#:764,314)(764,200)(720,200){1}
wire [11:0] w7;    //: /sn:0 {0}(#:357,83)(357,93)(352,93){1}
//: {2}(348,93)(#:252,93){3}
//: {4}(350,95)(350,155){5}
wire [11:0] IR_out;    //: /sn:0 {0}(#:208,555)(213,555){1}
//: {2}(214,555)(380,555)(380,498){3}
//: {4}(380,497)(380,490)(384,490)(384,469){5}
//: {6}(384,468)(384,436){7}
//: {8}(384,435)(384,404){9}
//: {10}(384,403)(384,359){11}
//: {12}(384,358)(384,307)(350,307)(#:350,176){13}
wire [8:0] PC_1;    //: /sn:0 {0}(#:159,326)(159,462)(142,462){1}
wire [7:0] acc_out0;    //: /sn:0 {0}(#:699,200)(666,200)(666,383){1}
//: {2}(#:668,385)(782,385)(782,343){3}
//: {4}(666,387)(666,496){5}
wire w14;    //: /sn:0 {0}(108,325)(108,311)(135,311){1}
wire w4;    //: /sn:0 {0}(260,471)(189,471)(189,439)(126,439)(126,449){1}
wire w3;    //: /sn:0 {0}(331,471)(281,471){1}
wire [1:0] ALU_Ctrl_out;    //: /sn:0 {0}(#:482,402)(806,402)(806,327)(787,327){1}
wire [8:0] PC_input;    //: /sn:0 {0}(#:113,472)(20,472)(20,198)(59,198){1}
wire [4:0] ram_in;    //: /sn:0 {0}(388,359)(#:492,359)(492,82)(526,82){1}
wire [8:0] pcout;    //: /sn:0 {0}(#:143,297)(143,210)(124,210)(124,200){1}
//: {2}(126,198)(127,198)(127,131){3}
//: {4}(129,129)(139,129)(139,95)(#:217,95){5}
//: {6}(127,127)(127,121){7}
//: {8}(122,198)(#:80,198){9}
wire [8:0] IR_mx_IN;    //: /sn:0 {0}(#:214,550)(214,482)(142,482){1}
wire [7:0] w23;    //: /sn:0 {0}(#:770,358)(770,343){1}
wire [7:0] RAM_out;    //: /sn:0 {0}(#:561,80)(634,80)(634,496){1}
wire w22;    //: /sn:0 {0}(626,510)(611,510){1}
wire CLK;    //: /sn:0 {0}(279,217)(305,217)(305,194){1}
//: {2}(307,192)(515,192)(515,152)(710,152)(710,162){3}
//: {4}(305,190)(305,165)(313,165){5}
//: {6}(303,192)(224,192)(224,244){7}
//: {8}(222,246)(70,246)(70,236){9}
//: {10}(224,248)(224,261)(248,261){11}
wire [5:0] alu_ctrl_in;    //: /sn:0 {0}(#:388,404)(447,404){1}
wire w2;    //: /sn:0 {0}(375,498)(368,498)(368,505)(317,505)(317,476)(281,476){1}
wire w5;    //: /sn:0 {0}(281,466)(321,466)(321,451)(375,451)(375,436)(379,436){1}
wire [7:0] add_out;    //: /sn:0 {0}(#:650,525)(650,535)(746,535)(746,343){1}
//: enddecls

  _GGREG9 #(10, 10, 20) g8 (.Q(pcout), .D(PC_input), .EN(w0), .CLR(w13), .CK(CLK));   //: @(70,198) /sn:0 /R:1 /w:[ 9 1 5 1 9 ]
  //: VDD g4 (w8) @(456,135) /sn:0 /w:[ 5 ]
  //: SWITCH g13 (w0) @(29,48) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGREG12 #(10, 10, 20) g3 (.Q(IR_out), .D(w7), .EN(w11), .CLR(w8), .CK(CLK));   //: @(350,165) /sn:0 /w:[ 13 5 7 0 5 ]
  //: comment g34 @(723,172) /sn:0
  //: /line:"Working register (accumulator)"
  //: /end
  _GGADD8 #(68, 70, 62, 64) g37 (.A(RAM_out), .B(acc_out0), .S(add_out), .CI(w18), .CO(w22));   //: @(650,512) /sn:0 /w:[ 1 5 0 5 0 ]
  //: joint g51 (w18) @(689, 317) /w:[ 2 1 -1 4 ]
  //: SWITCH g2 (w1) @(212,160) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g1 (w7) @(350, 93) /w:[ 1 -1 2 4 ]
  //: joint g11 (CLK) @(305, 192) /w:[ 2 4 6 1 ]
  //: comment g16 @(358,176) /sn:0
  //: /line:"Instruction register"
  //: /line:""
  //: /end
  //: LED g28 (CLK) @(255,261) /sn:0 /R:3 /w:[ 11 ] /type:0
  //: joint g10 (pcout) @(127, 129) /w:[ 4 6 -1 3 ]
  //: GROUND g50 (w18) @(689,296) /sn:0 /R:2 /w:[ 0 ]
  assign w2 = IR_out[9]; //: TAP g32 @(378,498) /sn:0 /R:2 /w:[ 0 3 4 ] /ss:0
  _GGAND3 #(8) g19 (.I0(w2), .I1(w3), .I2(w5), .Z(w4));   //: @(270,471) /sn:0 /R:2 /w:[ 1 1 0 0 ]
  //: joint g27 (w9) @(175, 290) /w:[ 1 2 -1 4 ]
  _GGRAM5x8 #(10, 60, 70, 10, 10, 10) g38 (.A(ram_in), .D(RAM_out), .WE(w8), .OE(w11), .CS(w11));   //: @(544,81) /sn:0 /w:[ 1 0 3 11 13 ]
  _GGCLOCK_P100_0_50 g6 (.Z(CLK));   //: @(266,217) /sn:0 /w:[ 0 ] /omega:100 /phi:0 /duty:50
  //: DIP g53 (w10) @(882,617) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g9 (w7) @(357,76) /sn:0 /w:[ 0 ] /type:1
  assign IR_mx_IN = IR_out[9:0]; //: TAP g7 @(214,553) /sn:0 /R:1 /w:[ 0 1 2 ] /ss:0
  assign w6 = IR_out[10]; //: TAP g31 @(382,469) /sn:0 /R:2 /w:[ 0 5 6 ] /ss:0
  //: joint g20 (pcout) @(124, 198) /w:[ 2 -1 8 1 ]
  //: comment g15 @(192,52) /sn:0
  //: /line:"Program memory"
  //: /end
  assign ram_in = IR_out[4:0]; //: TAP g39 @(382,359) /sn:0 /R:2 /w:[ 0 11 12 ] /ss:1
  //: joint g43 (w8) @(445, 155) /w:[ 2 4 -1 1 ]
  //: comment g48 @(434,364) /sn:0
  //: /line:"ALU Control"
  //: /end
  _GGNBUF #(2) g25 (.I(w6), .Z(w3));   //: @(341,471) /sn:0 /R:2 /w:[ 1 0 ]
  //: joint g29 (CLK) @(224, 246) /w:[ -1 7 8 10 ]
  _GGADD9 #(76, 78, 70, 72) g17 (.A(pcout), .B(w9), .S(PC_1), .CI(w16), .CO(w14));   //: @(159,313) /sn:0 /w:[ 0 5 0 1 1 ]
  //: joint g42 (w11) @(537, 121) /w:[ 10 12 9 -1 ]
  //: VDD g52 (w15) @(745,224) /sn:0 /w:[ 0 ]
  //: GROUND g5 (w11) @(445,91) /sn:0 /R:1 /w:[ 0 ]
  //: comment g14 @(95,208) /sn:0
  //: /line:"Program counter"
  //: /line:""
  //: /end
  _GGMUX4x8 #(12, 12) g44 (.I0(acc_out0), .I1(w23), .I2(w10), .I3(add_out), .S(ALU_Ctrl_out), .Z(acc_in));   //: @(764,327) /sn:0 /R:2 /w:[ 3 1 1 1 1 0 ] /ss:0 /do:0
  //: joint g47 (w11) @(402, 170) /w:[ 4 3 6 -1 ]
  //: joint g24 (w0) @(98, 48) /w:[ 2 -1 1 4 ]
  //: SWITCH g21 (w13) @(30,94) /sn:0 /w:[ 0 ] /st:1 /dn:1
  //: comment g36 @(527,257) /sn:0
  //: /line:"ALU"
  //: /end
  //: LED g23 (w0) @(130,15) /sn:0 /w:[ 3 ] /type:0
  //: joint g41 (w11) @(420, 91) /w:[ 1 -1 2 8 ]
  //: comment g40 @(563,39) /sn:0
  //: /line:"File register (RAM)"
  //: /end
  //: LED g26 (w14) @(108,332) /sn:0 /R:2 /w:[ 0 ] /type:0
  //: GROUND g22 (w16) @(206,336) /sn:0 /w:[ 0 ]
  _GGROM9x12 #(10, 30) g0 (.A(pcout), .D(w7), .OE(w1));   //: @(235,94) /sn:0 /w:[ 5 3 1 ] /mem:"/home/lelu0/oiakp/program.mem"
  //: frame g35 @(527,275) /sn:0 /wi:544 /ht:307 /tx:""
  _GGROM6x2 #(10, 30) g45 (.A(alu_ctrl_in), .D(ALU_Ctrl_out), .OE(w11));   //: @(465,403) /sn:0 /w:[ 1 0 5 ] /mem:"/home/lelu0/oiakp/alucntrl.mem"
  assign alu_ctrl_in = IR_out[11:6]; //: TAP g46 @(382,404) /sn:0 /R:2 /w:[ 0 9 10 ] /ss:1
  //: DIP g18 (w9) @(317,372) /sn:0 /R:2 /w:[ 0 ] /st:1 /dn:1
  _GGMUX2x9 #(8, 8) g12 (.I0(PC_1), .I1(IR_mx_IN), .S(w4), .Z(PC_input));   //: @(126,472) /sn:0 /R:3 /w:[ 1 1 1 0 ] /ss:0 /do:0
  assign w5 = IR_out[11]; //: TAP g30 @(382,436) /sn:0 /R:2 /w:[ 1 7 8 ] /ss:0
  _GGREG8 #(10, 10, 20) g33 (.Q(acc_out0), .D(acc_in), .EN(w18), .CLR(w15), .CK(CLK));   //: @(710,200) /sn:0 /R:3 /w:[ 0 1 3 1 3 ]
  //: joint g49 (acc_out0) @(666, 385) /w:[ 2 1 -1 4 ]

endmodule
//: /netlistEnd

//: /netlistBegin ROM
module ROM();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
reg [7:0] w1;    //: /sn:0 {0}(#:92,155)(92,159){1}
//: {2}(94,161)(#:104,161)(104,250)(169,250){3}
//: {4}(92,163)(92,172){5}
reg w2;    //: /sn:0 {0}(121,324)(175,324)(175,282)(185,282){1}
//: {2}(187,280)(187,275){3}
//: {4}(187,284)(187,292){5}
wire [7:0] w0;    //: /sn:0 {0}(#:204,248)(267,248)(267,166)(277,166){1}
//: {2}(279,164)(279,158){3}
//: {4}(279,168)(#:279,175){5}
//: enddecls

  //: joint g4 (w0) @(279, 166) /w:[ -1 2 1 4 ]
  //: joint g3 (w1) @(92, 161) /w:[ 2 1 -1 4 ]
  _GGROM8x8 #(10, 30) g2 (.A(w1), .D(w0), .OE(w2));   //: @(187,249) /sn:0 /w:[ 3 0 3 ]
  //: DIP g1 (w1) @(92,145) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g6 (w2) @(187, 282) /w:[ -1 2 1 4 ]
  //: SWITCH g5 (w2) @(104,324) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g0 (w0) @(279,151) /sn:0 /w:[ 3 ] /type:1

endmodule
//: /netlistEnd

