//: version "2.0-b10"
//: property encoding = "iso8859-1"
//: property locale = "en"
//: property prefix = "_GG"
//: property title = "pic.v"
//: property timingViolationMode = 2
//: property initTime = "0 ns"

`timescale 1ns/1ns

//: /netlistBegin main
module main;    //: root_module
reg [1:0] w32;    //: /sn:0 {0}(#:1037,361)(1037,415)(969,415)(969,424){1}
reg [7:0] w7;    //: /sn:0 {0}(776,358)(776,679)(1000,679)(#:1000,632){1}
supply0 w16;    //: /sn:0 {0}(206,330)(206,311)(183,311){1}
supply1 w15;    //: /sn:0 {0}(715,238)(715,248)(734,248)(734,224){1}
supply0 w0;    //: /sn:0 {0}(101,150)(101,145)(75,145)(75,160){1}
reg w1;    //: /sn:0 {0}(229,160)(235,160)(235,120){1}
supply0 w18;    //: /sn:0 {0}(674,510)(689,510)(689,476){1}
//: {2}(689,472)(689,315){3}
//: {4}(689,311)(689,302){5}
//: {6}(687,313)(595,313)(595,323){7}
//: {8}(687,474)(583,474)(583,439){9}
supply1 w8;    //: /sn:0 {0}(585,323)(585,298)(595,298)(595,139)(479,139){1}
//: {2}(477,137)(477,45)(544,45)(544,57){3}
//: {4}(477,141)(477,155)(447,155){5}
//: {6}(445,153)(445,135){7}
//: {8}(445,157)(445,160)(389,160){9}
supply0 w11;    //: /sn:0 {0}(466,429)(466,441)(420,441)(420,170)(404,170){1}
//: {2}(402,168)(402,91)(418,91){3}
//: {4}(422,91)(439,91){5}
//: {6}(420,93)(420,121)(535,121){7}
//: {8}(539,121)(551,121)(551,107){9}
//: {10}(537,119)(537,107){11}
//: {12}(400,170)(389,170){13}
reg [7:0] w10;    //: /sn:0 {0}(770,358)(770,646)(882,646)(#:882,627){1}
reg w13;    //: /sn:0 {0}(47,94)(53,94){1}
//: {2}(57,94)(65,94)(65,160){3}
//: {4}(55,96)(55,643)(606,643)(606,423)(596,423){5}
reg [8:0] w9;    //: /sn:0 {0}(#:317,361)(317,290)(177,290){1}
//: {2}(175,288)(#:175,283){3}
//: {4}(175,292)(175,297){5}
wire [7:0] acc_in;    //: /sn:0 {0}(#:862,167)(862,155)(771,155)(771,182){1}
//: {2}(#:769,184)(727,184)(727,395)(783,395)(783,358){3}
//: {4}(771,186)(771,200)(720,200){5}
wire w6;    //: /sn:0 {0}(379,469)(372,469)(372,471)(347,471){1}
wire [8:0] PC_1;    //: /sn:0 {0}(#:159,326)(159,462)(142,462){1}
wire [11:0] IR_out;    //: /sn:0 {0}(#:1195,9)(1195,12)(959,12){1}
//: {2}(958,12)(920,12){3}
//: {4}(919,12)(894,12){5}
//: {6}(893,12)(869,12){7}
//: {8}(868,12)(835,12){9}
//: {10}(834,12)(281,12)(281,212)(#:348,212){11}
//: {12}(350,210)(#:350,176){13}
//: {14}(350,214)(350,320)(384,320)(384,358){15}
//: {16}(384,359)(384,404){17}
//: {18}(384,405)(384,435){19}
//: {20}(384,436)(384,468){21}
//: {22}(384,469)(384,497){23}
//: {24}(384,498)(384,525){25}
//: {26}(384,526)(384,541){27}
//: {28}(384,542)(384,555)(372,555){29}
//: {30}(371,555)(350,555){31}
//: {32}(349,555)(294,555){33}
//: {34}(293,555)(214,555){35}
//: {36}(213,555)(#:208,555){37}
wire w45;    //: /sn:0 {0}(920,16)(920,24)(912,24)(912,105){1}
wire w14;    //: /sn:0 {0}(108,325)(108,311)(135,311){1}
wire w19;    //: /sn:0 {0}(70,236)(70,246)(224,246)(224,192)(303,192){1}
//: {2}(307,192)(513,192){3}
//: {4}(517,192)(549,192)(549,358)(590,358)(590,355){5}
//: {6}(515,190)(515,150)(710,150)(710,162){7}
//: {8}(305,190)(305,165)(313,165){9}
//: {10}(305,194)(305,217)(279,217){11}
wire w4;    //: /sn:0 {0}(260,471)(189,471)(189,439)(126,439)(126,449){1}
wire [7:0] w38;    //: /sn:0 {0}(#:750,373)(750,358){1}
wire [7:0] w51;    //: /sn:0 {0}(#:964,430)(964,456)(875,456)(#:875,424){1}
wire w3;    //: /sn:0 {0}(331,471)(281,471){1}
wire xor_mux_cntrl;    //: /sn:0 {0}(905,126)(905,180)(885,180){1}
wire [7:0] w37;    //: /sn:0 {0}(#:756,373)(756,358){1}
wire [7:0] w34;    //: /sn:0 {0}(#:800,261)(800,297)(832,297)(832,575)(#:294,575)(294,559){1}
wire [8:0] PC_input;    //: /sn:0 {0}(#:113,472)(20,472)(20,198)(59,198){1}
wire [7:0] w43;    //: /sn:0 {0}(870,424)(870,456)(#:668,456){1}
//: {2}(666,454)(#:666,261){3}
//: {4}(666,458)(#:666,496){5}
wire [4:0] ram_in;    //: /sn:0 {0}(388,359)(#:492,359)(492,82)(526,82){1}
wire [7:0] w31;    //: /sn:0 {0}(#:760,329)(760,306)(820,306)(820,261){1}
wire W_write_ctrl;    //: /sn:0 {0}(606,334)(705,334)(705,238){1}
wire w28;    //: /sn:0 {0}(438,537)(372,537)(372,550){1}
wire [7:0] movlw_mux_out;    //: /sn:0 {0}(852,196)(852,228)(#:810,228)(#:810,232){1}
wire w24;    //: /sn:0 {0}(350,550)(350,532)(438,532){1}
wire w23;    //: /sn:0 {0}(388,526)(396,526)(396,527)(438,527){1}
wire [8:0] IR_mx_IN;    //: /sn:0 {0}(#:214,550)(214,482)(142,482){1}
wire [8:0] pcout;    //: /sn:0 {0}(#:143,297)(143,210)(124,210)(124,200){1}
//: {2}(126,198)(127,198)(127,131){3}
//: {4}(129,129)(139,129)(139,95)(#:217,95){5}
//: {6}(127,127)(127,121){7}
//: {8}(122,198)(#:80,198){9}
wire [7:0] w36;    //: /sn:0 {0}(763,358)(763,534)(650,534)(#:650,525){1}
wire [2:0] w41;    //: /sn:0 {0}(#:483,402)(813,402)(813,342)(783,342){1}
wire w20;    //: /sn:0 {0}(606,344)(616,344)(616,449)(563,449)(563,439){1}
wire [7:0] RAM_out;    //: /sn:0 {0}(#:561,80)(634,80)(634,496){1}
wire [7:0] w40;    //: /sn:0 {0}(#:736,373)(736,358){1}
wire w30;    //: /sn:0 {0}(438,542)(388,542){1}
wire w22;    //: /sn:0 {0}(626,510)(611,510){1}
wire w17;    //: /sn:0 {0}(573,410)(573,369)(564,369)(564,339)(574,339){1}
wire [5:0] alu_ctrl_in;    //: /sn:0 {0}(#:388,405)(418,405)(418,404)(448,404){1}
wire [5:0] ir_xor_pipe;    //: /sn:0 {0}(#:959,16)(959,424){1}
wire w2;    //: /sn:0 {0}(379,498)(372,498)(372,505)(321,505)(321,476)(281,476){1}
wire w49;    //: /sn:0 {0}(902,105)(902,40)(869,40)(869,16){1}
wire w27;    //: /sn:0 {0}(459,534)(568,534)(568,564)(848,564)(848,245)(833,245){1}
wire w5;    //: /sn:0 {0}(281,466)(321,466)(321,451)(375,451)(375,436)(379,436){1}
wire [7:0] acc_out;    //: /sn:0 {0}(#:699,200)(666,200)(666,245){1}
wire [11:0] Program;    //: /sn:0 {0}(#:357,83)(357,93)(352,93){1}
//: {2}(348,93)(#:252,93){3}
//: {4}(350,95)(350,155){5}
wire w47;    //: /sn:0 {0}(894,16)(894,32)(907,32)(907,105){1}
wire w50;    //: /sn:0 {0}(897,105)(897,54)(835,54)(835,16){1}
wire [7:0] xor_out;    //: /sn:0 {0}(872,196)(#:872,403){1}
wire [7:0] w39;    //: /sn:0 {0}(#:743,373)(743,358){1}
//: enddecls

  //: LED g61 (IR_out) @(1195,2) /sn:0 /w:[ 0 ] /type:1
  //: VDD g4 (w8) @(456,135) /sn:0 /w:[ 7 ]
  _GGREG9 #(10, 10, 20) g8 (.Q(pcout), .D(PC_input), .EN(w0), .CLR(w13), .CK(w19));   //: @(70,198) /sn:0 /R:1 /w:[ 9 1 1 3 0 ]
  //: GROUND g13 (w0) @(101,156) /sn:0 /w:[ 0 ]
  _GGADD8 #(68, 70, 62, 64) g37 (.A(RAM_out), .B(w43), .S(w36), .CI(w18), .CO(w22));   //: @(650,512) /sn:0 /w:[ 1 5 1 0 0 ]
  //: comment g34 @(643,129) /sn:0
  //: /line:"Working register (accumulator)"
  //: /end
  _GGREG12 #(10, 10, 20) g3 (.Q(IR_out), .D(Program), .EN(w11), .CLR(w8), .CK(w19));   //: @(350,165) /sn:0 /w:[ 13 5 13 9 9 ]
  //: joint g51 (w19) @(515, 192) /w:[ 4 6 3 -1 ]
  //: joint g55 (w8) @(477, 139) /w:[ 1 2 -1 4 ]
  //: joint g58 (w13) @(55, 94) /w:[ 2 -1 1 4 ]
  assign w30 = IR_out[11]; //: TAP g65 @(382,542) /sn:0 /R:2 /w:[ 1 28 27 ] /ss:1
  //: SWITCH g2 (w1) @(212,160) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g76 (acc_in) @(771, 184) /w:[ -1 1 2 4 ]
  //: joint g59 (w18) @(689, 474) /w:[ -1 2 8 1 ]
  //: joint g1 (Program) @(350, 93) /w:[ 1 -1 2 4 ]
  //: joint g72 (w43) @(666, 456) /w:[ 1 2 -1 4 ]
  _GGNOR4 #(10) g64 (.I0(w23), .I1(w24), .I2(!w28), .I3(!w30), .Z(w27));   //: @(449,534) /sn:0 /w:[ 1 1 0 0 0 ]
  //: comment g16 @(358,176) /sn:0
  //: /line:"Instruction register"
  //: /line:""
  //: /end
  //: joint g11 (w19) @(305, 192) /w:[ 2 8 1 10 ]
  //: GROUND g50 (w18) @(689,296) /sn:0 /R:2 /w:[ 5 ]
  //: joint g10 (pcout) @(127, 129) /w:[ 4 6 -1 3 ]
  assign w51 = {w32, ir_xor_pipe}; //: CONCAT g78  @(964,429) /sn:0 /R:3 /w:[ 0 1 1 ] /dr:0 /tp:0 /drp:1
  //: joint g27 (w9) @(175, 290) /w:[ 1 2 -1 4 ]
  _GGAND3 #(8) g19 (.I0(w2), .I1(w3), .I2(w5), .Z(w4));   //: @(270,471) /sn:0 /R:2 /w:[ 1 1 0 0 ]
  assign w2 = IR_out[9]; //: TAP g32 @(382,498) /sn:0 /R:2 /w:[ 0 24 23 ] /ss:0
  _GGMUX2x8 #(8, 8) g69 (.I0(w31), .I1(w34), .S(w27), .Z(movlw_mux_out));   //: @(810,245) /sn:0 /R:2 /w:[ 1 0 1 1 ] /ss:0 /do:0
  _GGCLOCK_P100_0_50 g6 (.Z(w19));   //: @(266,217) /sn:0 /w:[ 11 ] /omega:100 /phi:0 /duty:50
  _GGRAM5x8 #(10, 60, 70, 10, 10, 10) g38 (.A(ram_in), .D(RAM_out), .WE(w8), .OE(w11), .CS(w11));   //: @(544,81) /sn:0 /w:[ 1 0 3 9 11 ]
  assign IR_mx_IN = IR_out[9:0]; //: TAP g7 @(214,553) /sn:0 /R:1 /w:[ 0 36 35 ] /ss:0
  //: LED g9 (Program) @(357,76) /sn:0 /w:[ 0 ] /type:1
  //: DIP g53 (w10) @(882,617) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: DIP g75 (w32) @(1037,351) /sn:0 /w:[ 0 ] /st:0 /dn:1
  _GGMUX2 #(8, 8) g57 (.I0(w18), .I1(w20), .S(w13), .Z(w17));   //: @(573,423) /sn:0 /R:2 /w:[ 9 1 5 0 ] /ss:0 /do:0
  //: comment g15 @(192,52) /sn:0
  //: /line:"Program memory"
  //: /end
  //: joint g20 (pcout) @(124, 198) /w:[ 2 -1 8 1 ]
  assign w6 = IR_out[10]; //: TAP g31 @(382,469) /sn:0 /R:2 /w:[ 0 22 21 ] /ss:0
  _GGXOR2x8 #(8) g71 (.I0(w43), .I1(w51), .Z(xor_out));   //: @(872,413) /sn:0 /R:1 /w:[ 0 1 1 ]
  assign w24 = IR_out[9]; //: TAP g68 @(350,553) /sn:0 /R:1 /w:[ 0 32 31 ] /ss:0
  assign w28 = IR_out[10]; //: TAP g67 @(372,553) /sn:0 /R:1 /w:[ 1 30 29 ] /ss:0
  assign ram_in = IR_out[4:0]; //: TAP g39 @(382,359) /sn:0 /R:2 /w:[ 0 16 15 ] /ss:1
  //: comment g48 @(434,364) /sn:0
  //: /line:"ALU Control"
  //: /end
  //: joint g43 (w8) @(445, 155) /w:[ 5 6 -1 8 ]
  //: joint g62 (IR_out) @(350, 212) /w:[ -1 12 11 14 ]
  _GGADD9 #(76, 78, 70, 72) g17 (.A(pcout), .B(w9), .S(PC_1), .CI(w16), .CO(w14));   //: @(159,313) /sn:0 /w:[ 0 5 0 1 1 ]
  _GGNBUF #(2) g25 (.I(w6), .Z(w3));   //: @(341,471) /sn:0 /R:2 /w:[ 1 0 ]
  assign ir_xor_pipe = IR_out[5:0]; //: TAP g73 @(959,10) /sn:0 /R:1 /w:[ 0 2 1 ] /ss:1
  //: DIP g63 (w7) @(1000,622) /sn:0 /w:[ 1 ] /st:0 /dn:1
  //: VDD g52 (w15) @(745,224) /sn:0 /w:[ 1 ]
  //: joint g42 (w11) @(537, 121) /w:[ 8 10 7 -1 ]
  assign w49 = IR_out[9]; //: TAP g83 @(869,10) /sn:0 /R:1 /w:[ 1 8 7 ] /ss:1
  //: comment g14 @(95,208) /sn:0
  //: /line:"Program counter"
  //: /line:""
  //: /end
  //: GROUND g5 (w11) @(445,91) /sn:0 /R:1 /w:[ 5 ]
  //: joint g56 (w18) @(689, 313) /w:[ -1 4 6 3 ]
  //: joint g47 (w11) @(402, 170) /w:[ 1 2 12 -1 ]
  _GGMUX8x8 #(20, 20) g44 (.I0(acc_in), .I1(w7), .I2(w10), .I3(w36), .I4(w37), .I5(w38), .I6(w39), .I7(w40), .S(w41), .Z(w31));   //: @(760,342) /sn:0 /R:2 /w:[ 3 0 0 0 1 1 1 1 1 0 ] /ss:0 /do:0
  _GGMUX2x8 #(8, 8) g79 (.I0(movlw_mux_out), .I1(xor_out), .S(xor_mux_cntrl), .Z(acc_in));   //: @(862,180) /sn:0 /R:2 /w:[ 0 0 1 0 ] /ss:0 /do:1
  _GGAND4 #(10) g80 (.I0(w45), .I1(w47), .I2(w49), .I3(w50), .Z(xor_mux_cntrl));   //: @(905,116) /sn:0 /R:3 /w:[ 1 1 0 0 0 ]
  //: comment g36 @(527,257) /sn:0
  //: /line:"ALU"
  //: /end
  //: SWITCH g21 (w13) @(30,94) /sn:0 /w:[ 0 ] /st:1 /dn:1
  assign w50 = IR_out[8]; //: TAP g84 @(835,10) /sn:0 /R:1 /w:[ 1 10 9 ] /ss:1
  //: joint g41 (w11) @(420, 91) /w:[ 4 -1 3 6 ]
  //: comment g40 @(563,39) /sn:0
  //: /line:"File register (RAM)"
  //: /end
  assign w45 = IR_out[11]; //: TAP g81 @(920,10) /sn:0 /R:1 /w:[ 0 4 3 ] /ss:1
  _GGBUF8 #(4) g60 (.I(acc_out), .Z(w43));   //: @(666,251) /sn:0 /R:3 /w:[ 1 3 ]
  _GGFF #(10, 10, 20) g54 (.Q(W_write_ctrl), ._Q(w20), .D(w17), .EN(w18), .CLR(w8), .CK(w19));   //: @(590,339) /sn:0 /w:[ 0 0 1 7 0 5 ] /mi:0
  assign w34 = IR_out[7:0]; //: TAP g70 @(294,553) /sn:0 /R:1 /w:[ 1 34 33 ] /ss:1
  assign alu_ctrl_in = IR_out[11:6]; //: TAP g46 @(382,405) /sn:0 /R:2 /w:[ 0 18 17 ] /ss:1
  _GGROM6x3 #(10, 30) g45 (.A(alu_ctrl_in), .D(w41), .OE(w11));   //: @(466,403) /sn:0 /w:[ 1 0 0 ] /mem:"/home/lelu0/oiakp/alucntrl.mem"
  //: frame g35 @(533,275) /sn:0 /wi:544 /ht:307 /tx:""
  _GGROM9x12 #(10, 30) g0 (.A(pcout), .D(Program), .OE(w1));   //: @(235,94) /sn:0 /w:[ 5 3 1 ] /mem:"/home/lelu0/oiakp/program.mem"
  //: GROUND g22 (w16) @(206,336) /sn:0 /w:[ 0 ]
  //: LED g26 (w14) @(108,332) /sn:0 /R:2 /w:[ 0 ] /type:0
  assign w23 = IR_out[8]; //: TAP g66 @(382,526) /sn:0 /R:2 /w:[ 0 26 25 ] /ss:1
  assign w47 = IR_out[10]; //: TAP g82 @(894,10) /sn:0 /R:1 /w:[ 0 6 5 ] /ss:1
  _GGMUX2x9 #(8, 8) g12 (.I0(PC_1), .I1(IR_mx_IN), .S(w4), .Z(PC_input));   //: @(126,472) /sn:0 /R:3 /w:[ 1 1 1 0 ] /ss:0 /do:0
  //: DIP g18 (w9) @(317,372) /sn:0 /R:2 /w:[ 0 ] /st:1 /dn:1
  _GGREG8 #(20, 20, 40) g33 (.Q(acc_out), .D(acc_in), .EN(W_write_ctrl), .CLR(w15), .CK(w19));   //: @(710,200) /sn:0 /R:3 /delay:" 20 20 40" /w:[ 0 5 1 0 7 ]
  assign w5 = IR_out[11]; //: TAP g30 @(382,436) /sn:0 /R:2 /w:[ 1 20 19 ] /ss:0
  //: comment g49 @(973,589) /sn:0
  //: /line:"const. zero"
  //: /end

endmodule
//: /netlistEnd

//: /netlistBegin ROM
module ROM();
//: interface  /sz:(40, 40) /bd:[ ] /pd: 0 /pi: 0 /pe: 1 /pp: 1
reg [7:0] w1;    //: /sn:0 {0}(#:92,155)(92,159){1}
//: {2}(94,161)(#:104,161)(104,250)(169,250){3}
//: {4}(92,163)(92,172){5}
reg w2;    //: /sn:0 {0}(121,324)(175,324)(175,282)(185,282){1}
//: {2}(187,280)(187,275){3}
//: {4}(187,284)(187,292){5}
wire [7:0] w0;    //: /sn:0 {0}(#:204,248)(267,248)(267,166)(277,166){1}
//: {2}(279,164)(279,158){3}
//: {4}(279,168)(#:279,175){5}
//: enddecls

  //: joint g4 (w0) @(279, 166) /w:[ -1 2 1 4 ]
  //: joint g3 (w1) @(92, 161) /w:[ 2 1 -1 4 ]
  _GGROM8x8 #(10, 30) g2 (.A(w1), .D(w0), .OE(w2));   //: @(187,249) /sn:0 /w:[ 3 0 3 ]
  //: DIP g1 (w1) @(92,145) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: joint g6 (w2) @(187, 282) /w:[ -1 2 1 4 ]
  //: SWITCH g5 (w2) @(104,324) /sn:0 /w:[ 0 ] /st:0 /dn:1
  //: LED g0 (w0) @(279,151) /sn:0 /w:[ 3 ] /type:1

endmodule
//: /netlistEnd

